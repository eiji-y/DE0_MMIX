// MMIX_system.v

// Generated using ACDS version 13.1 182 at 2017.12.13.20:05:13

`timescale 1 ps / 1 ps
module MMIX_system (
		input  wire        clk_clk,          //        clk.clk
		input  wire        reset_reset_n,    //      reset.reset_n
		output wire [11:0] sdram_wire_addr,  // sdram_wire.addr
		output wire [1:0]  sdram_wire_ba,    //           .ba
		output wire        sdram_wire_cas_n, //           .cas_n
		output wire        sdram_wire_cke,   //           .cke
		output wire        sdram_wire_cs_n,  //           .cs_n
		inout  wire [15:0] sdram_wire_dq,    //           .dq
		output wire [1:0]  sdram_wire_dqm,   //           .dqm
		output wire        sdram_wire_ras_n, //           .ras_n
		output wire        sdram_wire_we_n,  //           .we_n
		output wire        sdram_clk_clk,    //  sdram_clk.clk
		output wire [31:0] dbg_led_led,      //    dbg_led.led
		input  wire        dbg_led_btn,      //           .btn
		output wire [21:0] flash_wire_ADDR,  // flash_wire.ADDR
		output wire        flash_wire_CE_N,  //           .CE_N
		output wire        flash_wire_OE_N,  //           .OE_N
		output wire        flash_wire_WE_N,  //           .WE_N
		output wire        flash_wire_RST_N, //           .RST_N
		inout  wire [7:0]  flash_wire_DQ,    //           .DQ
		output wire        vga_wire_CLK,     //   vga_wire.CLK
		output wire        vga_wire_HS,      //           .HS
		output wire        vga_wire_VS,      //           .VS
		output wire [3:0]  vga_wire_R,       //           .R
		output wire [3:0]  vga_wire_G,       //           .G
		output wire [3:0]  vga_wire_B        //           .B
	);

	wire         clocks_sys_clk_clk;                                                                                  // clocks:sys_clk_clk -> [Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0:i_clock, mm_interconnect_0:clocks_sys_clk_clk, mmix_qsys_0:clk, rst_controller:clk, sdram:clk, video_character_buffer_with_dma_0:clk, video_dual_clock_buffer_0:clk_stream_in, video_pll_0:ref_clk_clk]
	wire         video_character_buffer_with_dma_0_avalon_char_source_endofpacket;                                    // video_character_buffer_with_dma_0:stream_endofpacket -> video_dual_clock_buffer_0:stream_in_endofpacket
	wire         video_character_buffer_with_dma_0_avalon_char_source_valid;                                          // video_character_buffer_with_dma_0:stream_valid -> video_dual_clock_buffer_0:stream_in_valid
	wire         video_character_buffer_with_dma_0_avalon_char_source_startofpacket;                                  // video_character_buffer_with_dma_0:stream_startofpacket -> video_dual_clock_buffer_0:stream_in_startofpacket
	wire  [29:0] video_character_buffer_with_dma_0_avalon_char_source_data;                                           // video_character_buffer_with_dma_0:stream_data -> video_dual_clock_buffer_0:stream_in_data
	wire         video_character_buffer_with_dma_0_avalon_char_source_ready;                                          // video_dual_clock_buffer_0:stream_in_ready -> video_character_buffer_with_dma_0:stream_ready
	wire         video_dual_clock_buffer_0_avalon_dc_buffer_source_endofpacket;                                       // video_dual_clock_buffer_0:stream_out_endofpacket -> video_vga_controller_0:endofpacket
	wire         video_dual_clock_buffer_0_avalon_dc_buffer_source_valid;                                             // video_dual_clock_buffer_0:stream_out_valid -> video_vga_controller_0:valid
	wire         video_dual_clock_buffer_0_avalon_dc_buffer_source_startofpacket;                                     // video_dual_clock_buffer_0:stream_out_startofpacket -> video_vga_controller_0:startofpacket
	wire  [29:0] video_dual_clock_buffer_0_avalon_dc_buffer_source_data;                                              // video_dual_clock_buffer_0:stream_out_data -> video_vga_controller_0:data
	wire         video_dual_clock_buffer_0_avalon_dc_buffer_source_ready;                                             // video_vga_controller_0:ready -> video_dual_clock_buffer_0:stream_out_ready
	wire         video_pll_0_vga_clk_clk;                                                                             // video_pll_0:vga_clk_clk -> [rst_controller_002:clk, video_dual_clock_buffer_0:clk_stream_out, video_vga_controller_0:clk]
	wire         mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_buffer_slave_waitrequest;            // video_character_buffer_with_dma_0:buf_waitrequest -> mm_interconnect_0:video_character_buffer_with_dma_0_avalon_char_buffer_slave_waitrequest
	wire   [7:0] mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_buffer_slave_writedata;              // mm_interconnect_0:video_character_buffer_with_dma_0_avalon_char_buffer_slave_writedata -> video_character_buffer_with_dma_0:buf_writedata
	wire  [12:0] mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_buffer_slave_address;                // mm_interconnect_0:video_character_buffer_with_dma_0_avalon_char_buffer_slave_address -> video_character_buffer_with_dma_0:buf_address
	wire         mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_buffer_slave_chipselect;             // mm_interconnect_0:video_character_buffer_with_dma_0_avalon_char_buffer_slave_chipselect -> video_character_buffer_with_dma_0:buf_chipselect
	wire         mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_buffer_slave_write;                  // mm_interconnect_0:video_character_buffer_with_dma_0_avalon_char_buffer_slave_write -> video_character_buffer_with_dma_0:buf_write
	wire         mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_buffer_slave_read;                   // mm_interconnect_0:video_character_buffer_with_dma_0_avalon_char_buffer_slave_read -> video_character_buffer_with_dma_0:buf_read
	wire   [7:0] mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_buffer_slave_readdata;               // video_character_buffer_with_dma_0:buf_readdata -> mm_interconnect_0:video_character_buffer_with_dma_0_avalon_char_buffer_slave_readdata
	wire   [0:0] mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_buffer_slave_byteenable;             // mm_interconnect_0:video_character_buffer_with_dma_0_avalon_char_buffer_slave_byteenable -> video_character_buffer_with_dma_0:buf_byteenable
	wire         mmix_qsys_0_master_waitrequest;                                                                      // mm_interconnect_0:mmix_qsys_0_master_waitrequest -> mmix_qsys_0:d_waitrequest
	wire  [63:0] mmix_qsys_0_master_writedata;                                                                        // mmix_qsys_0:d_writedata -> mm_interconnect_0:mmix_qsys_0_master_writedata
	wire  [27:0] mmix_qsys_0_master_address;                                                                          // mmix_qsys_0:d_address -> mm_interconnect_0:mmix_qsys_0_master_address
	wire         mmix_qsys_0_master_write;                                                                            // mmix_qsys_0:d_write -> mm_interconnect_0:mmix_qsys_0_master_write
	wire         mmix_qsys_0_master_read;                                                                             // mmix_qsys_0:d_read -> mm_interconnect_0:mmix_qsys_0_master_read
	wire  [63:0] mmix_qsys_0_master_readdata;                                                                         // mm_interconnect_0:mmix_qsys_0_master_readdata -> mmix_qsys_0:d_readdata
	wire         mmix_qsys_0_master_readdatavalid;                                                                    // mm_interconnect_0:mmix_qsys_0_master_readdatavalid -> mmix_qsys_0:d_readdatavalid
	wire   [7:0] mmix_qsys_0_master_byteenable;                                                                       // mmix_qsys_0:d_byteenable -> mm_interconnect_0:mmix_qsys_0_master_byteenable
	wire  [31:0] mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_control_slave_writedata;             // mm_interconnect_0:video_character_buffer_with_dma_0_avalon_char_control_slave_writedata -> video_character_buffer_with_dma_0:ctrl_writedata
	wire   [0:0] mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_control_slave_address;               // mm_interconnect_0:video_character_buffer_with_dma_0_avalon_char_control_slave_address -> video_character_buffer_with_dma_0:ctrl_address
	wire         mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_control_slave_chipselect;            // mm_interconnect_0:video_character_buffer_with_dma_0_avalon_char_control_slave_chipselect -> video_character_buffer_with_dma_0:ctrl_chipselect
	wire         mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_control_slave_write;                 // mm_interconnect_0:video_character_buffer_with_dma_0_avalon_char_control_slave_write -> video_character_buffer_with_dma_0:ctrl_write
	wire         mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_control_slave_read;                  // mm_interconnect_0:video_character_buffer_with_dma_0_avalon_char_control_slave_read -> video_character_buffer_with_dma_0:ctrl_read
	wire  [31:0] mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_control_slave_readdata;              // video_character_buffer_with_dma_0:ctrl_readdata -> mm_interconnect_0:video_character_buffer_with_dma_0_avalon_char_control_slave_readdata
	wire   [3:0] mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_control_slave_byteenable;            // mm_interconnect_0:video_character_buffer_with_dma_0_avalon_char_control_slave_byteenable -> video_character_buffer_with_dma_0:ctrl_byteenable
	wire         mm_interconnect_0_altera_up_flash_memory_ip_core_avalon_interface_0_flash_data_waitrequest;          // Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0:o_avalon_waitrequest -> mm_interconnect_0:Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_data_waitrequest
	wire  [31:0] mm_interconnect_0_altera_up_flash_memory_ip_core_avalon_interface_0_flash_data_writedata;            // mm_interconnect_0:Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_data_writedata -> Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0:i_avalon_writedata
	wire  [19:0] mm_interconnect_0_altera_up_flash_memory_ip_core_avalon_interface_0_flash_data_address;              // mm_interconnect_0:Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_data_address -> Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0:i_avalon_address
	wire         mm_interconnect_0_altera_up_flash_memory_ip_core_avalon_interface_0_flash_data_chipselect;           // mm_interconnect_0:Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_data_chipselect -> Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0:i_avalon_chip_select
	wire         mm_interconnect_0_altera_up_flash_memory_ip_core_avalon_interface_0_flash_data_write;                // mm_interconnect_0:Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_data_write -> Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0:i_avalon_write
	wire         mm_interconnect_0_altera_up_flash_memory_ip_core_avalon_interface_0_flash_data_read;                 // mm_interconnect_0:Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_data_read -> Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0:i_avalon_read
	wire  [31:0] mm_interconnect_0_altera_up_flash_memory_ip_core_avalon_interface_0_flash_data_readdata;             // Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0:o_avalon_readdata -> mm_interconnect_0:Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_data_readdata
	wire   [3:0] mm_interconnect_0_altera_up_flash_memory_ip_core_avalon_interface_0_flash_data_byteenable;           // mm_interconnect_0:Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_data_byteenable -> Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0:i_avalon_byteenable
	wire         mm_interconnect_0_sdram_s1_waitrequest;                                                              // sdram:za_waitrequest -> mm_interconnect_0:sdram_s1_waitrequest
	wire  [15:0] mm_interconnect_0_sdram_s1_writedata;                                                                // mm_interconnect_0:sdram_s1_writedata -> sdram:az_data
	wire  [21:0] mm_interconnect_0_sdram_s1_address;                                                                  // mm_interconnect_0:sdram_s1_address -> sdram:az_addr
	wire         mm_interconnect_0_sdram_s1_chipselect;                                                               // mm_interconnect_0:sdram_s1_chipselect -> sdram:az_cs
	wire         mm_interconnect_0_sdram_s1_write;                                                                    // mm_interconnect_0:sdram_s1_write -> sdram:az_wr_n
	wire         mm_interconnect_0_sdram_s1_read;                                                                     // mm_interconnect_0:sdram_s1_read -> sdram:az_rd_n
	wire  [15:0] mm_interconnect_0_sdram_s1_readdata;                                                                 // sdram:za_data -> mm_interconnect_0:sdram_s1_readdata
	wire         mm_interconnect_0_sdram_s1_readdatavalid;                                                            // sdram:za_valid -> mm_interconnect_0:sdram_s1_readdatavalid
	wire   [1:0] mm_interconnect_0_sdram_s1_byteenable;                                                               // mm_interconnect_0:sdram_s1_byteenable -> sdram:az_be_n
	wire         mm_interconnect_0_altera_up_flash_memory_ip_core_avalon_interface_0_flash_erase_control_waitrequest; // Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0:o_avalon_erase_waitrequest -> mm_interconnect_0:Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_erase_control_waitrequest
	wire  [31:0] mm_interconnect_0_altera_up_flash_memory_ip_core_avalon_interface_0_flash_erase_control_writedata;   // mm_interconnect_0:Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_erase_control_writedata -> Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0:i_avalon_erase_writedata
	wire         mm_interconnect_0_altera_up_flash_memory_ip_core_avalon_interface_0_flash_erase_control_chipselect;  // mm_interconnect_0:Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_erase_control_chipselect -> Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0:i_avalon_erase_chip_select
	wire         mm_interconnect_0_altera_up_flash_memory_ip_core_avalon_interface_0_flash_erase_control_write;       // mm_interconnect_0:Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_erase_control_write -> Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0:i_avalon_erase_write
	wire         mm_interconnect_0_altera_up_flash_memory_ip_core_avalon_interface_0_flash_erase_control_read;        // mm_interconnect_0:Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_erase_control_read -> Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0:i_avalon_erase_read
	wire  [31:0] mm_interconnect_0_altera_up_flash_memory_ip_core_avalon_interface_0_flash_erase_control_readdata;    // Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0:o_avalon_erase_readdata -> mm_interconnect_0:Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_erase_control_readdata
	wire   [3:0] mm_interconnect_0_altera_up_flash_memory_ip_core_avalon_interface_0_flash_erase_control_byteenable;  // mm_interconnect_0:Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_erase_control_byteenable -> Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0:i_avalon_erase_byteenable
	wire  [31:0] mmix_qsys_0_d_irq_irq;                                                                               // irq_mapper:sender_irq -> mmix_qsys_0:d_irq
	wire         rst_controller_reset_out_reset;                                                                      // rst_controller:reset_out -> [Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0:i_reset_n, mm_interconnect_0:mmix_qsys_0_reset_n_reset_bridge_in_reset_reset, mm_interconnect_0:sdram_reset_reset_bridge_in_reset_reset, sdram:reset_n, video_character_buffer_with_dma_0:reset, video_dual_clock_buffer_0:reset_stream_in, video_pll_0:ref_reset_reset]
	wire         rst_controller_001_reset_out_reset;                                                                  // rst_controller_001:reset_out -> clocks:ref_reset_reset
	wire         rst_controller_002_reset_out_reset;                                                                  // rst_controller_002:reset_out -> [video_dual_clock_buffer_0:reset_stream_out, video_vga_controller_0:reset]
	wire         video_pll_0_reset_source_reset;                                                                      // video_pll_0:reset_source_reset -> rst_controller_002:reset_in0

	mmix_qsys mmix_qsys_0 (
		.reset_n         (reset_reset_n),                    // reset_n.reset_n
		.clk             (clocks_sys_clk_clk),               //     clk.clk
		.d_irq           (mmix_qsys_0_d_irq_irq),            //   d_irq.irq
		.d_address       (mmix_qsys_0_master_address),       //  master.address
		.d_byteenable    (mmix_qsys_0_master_byteenable),    //        .byteenable
		.d_read          (mmix_qsys_0_master_read),          //        .read
		.d_readdata      (mmix_qsys_0_master_readdata),      //        .readdata
		.d_waitrequest   (mmix_qsys_0_master_waitrequest),   //        .waitrequest
		.d_write         (mmix_qsys_0_master_write),         //        .write
		.d_writedata     (mmix_qsys_0_master_writedata),     //        .writedata
		.d_readdatavalid (mmix_qsys_0_master_readdatavalid), //        .readdatavalid
		.dbg_led         (dbg_led_led),                      // conduit.export
		.dbg_btn         (dbg_led_btn)                       //        .export
	);

	MMIX_system_sdram sdram (
		.clk            (clocks_sys_clk_clk),                       //   clk.clk
		.reset_n        (~rst_controller_reset_out_reset),          // reset.reset_n
		.az_addr        (mm_interconnect_0_sdram_s1_address),       //    s1.address
		.az_be_n        (~mm_interconnect_0_sdram_s1_byteenable),   //      .byteenable_n
		.az_cs          (mm_interconnect_0_sdram_s1_chipselect),    //      .chipselect
		.az_data        (mm_interconnect_0_sdram_s1_writedata),     //      .writedata
		.az_rd_n        (~mm_interconnect_0_sdram_s1_read),         //      .read_n
		.az_wr_n        (~mm_interconnect_0_sdram_s1_write),        //      .write_n
		.za_data        (mm_interconnect_0_sdram_s1_readdata),      //      .readdata
		.za_valid       (mm_interconnect_0_sdram_s1_readdatavalid), //      .readdatavalid
		.za_waitrequest (mm_interconnect_0_sdram_s1_waitrequest),   //      .waitrequest
		.zs_addr        (sdram_wire_addr),                          //  wire.export
		.zs_ba          (sdram_wire_ba),                            //      .export
		.zs_cas_n       (sdram_wire_cas_n),                         //      .export
		.zs_cke         (sdram_wire_cke),                           //      .export
		.zs_cs_n        (sdram_wire_cs_n),                          //      .export
		.zs_dq          (sdram_wire_dq),                            //      .export
		.zs_dqm         (sdram_wire_dqm),                           //      .export
		.zs_ras_n       (sdram_wire_ras_n),                         //      .export
		.zs_we_n        (sdram_wire_we_n)                           //      .export
	);

	MMIX_system_clocks clocks (
		.ref_clk_clk        (clk_clk),                            //      ref_clk.clk
		.ref_reset_reset    (rst_controller_001_reset_out_reset), //    ref_reset.reset
		.sys_clk_clk        (clocks_sys_clk_clk),                 //      sys_clk.clk
		.sdram_clk_clk      (sdram_clk_clk),                      //    sdram_clk.clk
		.reset_source_reset ()                                    // reset_source.reset
	);

	Altera_UP_Flash_Memory_IP_Core_Avalon_Interface #(
		.FLASH_MEMORY_ADDRESS_WIDTH (22),
		.FLASH_MEMORY_WAIT_COUNT    (5)
	) altera_up_flash_memory_ip_core_avalon_interface_0 (
		.i_avalon_chip_select       (mm_interconnect_0_altera_up_flash_memory_ip_core_avalon_interface_0_flash_data_chipselect),           //          flash_data.chipselect
		.i_avalon_write             (mm_interconnect_0_altera_up_flash_memory_ip_core_avalon_interface_0_flash_data_write),                //                    .write
		.i_avalon_read              (mm_interconnect_0_altera_up_flash_memory_ip_core_avalon_interface_0_flash_data_read),                 //                    .read
		.i_avalon_address           (mm_interconnect_0_altera_up_flash_memory_ip_core_avalon_interface_0_flash_data_address),              //                    .address
		.i_avalon_byteenable        (mm_interconnect_0_altera_up_flash_memory_ip_core_avalon_interface_0_flash_data_byteenable),           //                    .byteenable
		.i_avalon_writedata         (mm_interconnect_0_altera_up_flash_memory_ip_core_avalon_interface_0_flash_data_writedata),            //                    .writedata
		.o_avalon_readdata          (mm_interconnect_0_altera_up_flash_memory_ip_core_avalon_interface_0_flash_data_readdata),             //                    .readdata
		.o_avalon_waitrequest       (mm_interconnect_0_altera_up_flash_memory_ip_core_avalon_interface_0_flash_data_waitrequest),          //                    .waitrequest
		.i_clock                    (clocks_sys_clk_clk),                                                                                  //          clock_sink.clk
		.i_reset_n                  (~rst_controller_reset_out_reset),                                                                     //    clock_sink_reset.reset_n
		.FL_ADDR                    (flash_wire_ADDR),                                                                                     //         conduit_end.export
		.FL_CE_N                    (flash_wire_CE_N),                                                                                     //                    .export
		.FL_OE_N                    (flash_wire_OE_N),                                                                                     //                    .export
		.FL_WE_N                    (flash_wire_WE_N),                                                                                     //                    .export
		.FL_RST_N                   (flash_wire_RST_N),                                                                                    //                    .export
		.FL_DQ                      (flash_wire_DQ),                                                                                       //                    .export
		.i_avalon_erase_write       (mm_interconnect_0_altera_up_flash_memory_ip_core_avalon_interface_0_flash_erase_control_write),       // flash_erase_control.write
		.i_avalon_erase_read        (mm_interconnect_0_altera_up_flash_memory_ip_core_avalon_interface_0_flash_erase_control_read),        //                    .read
		.i_avalon_erase_byteenable  (mm_interconnect_0_altera_up_flash_memory_ip_core_avalon_interface_0_flash_erase_control_byteenable),  //                    .byteenable
		.i_avalon_erase_writedata   (mm_interconnect_0_altera_up_flash_memory_ip_core_avalon_interface_0_flash_erase_control_writedata),   //                    .writedata
		.i_avalon_erase_chip_select (mm_interconnect_0_altera_up_flash_memory_ip_core_avalon_interface_0_flash_erase_control_chipselect),  //                    .chipselect
		.o_avalon_erase_readdata    (mm_interconnect_0_altera_up_flash_memory_ip_core_avalon_interface_0_flash_erase_control_readdata),    //                    .readdata
		.o_avalon_erase_waitrequest (mm_interconnect_0_altera_up_flash_memory_ip_core_avalon_interface_0_flash_erase_control_waitrequest)  //                    .waitrequest
	);

	MMIX_system_video_character_buffer_with_dma_0 video_character_buffer_with_dma_0 (
		.clk                  (clocks_sys_clk_clk),                                                                       //               clock_reset.clk
		.reset                (rst_controller_reset_out_reset),                                                           //         clock_reset_reset.reset
		.ctrl_address         (mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_control_slave_address),    // avalon_char_control_slave.address
		.ctrl_byteenable      (mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_control_slave_byteenable), //                          .byteenable
		.ctrl_chipselect      (mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_control_slave_chipselect), //                          .chipselect
		.ctrl_read            (mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_control_slave_read),       //                          .read
		.ctrl_write           (mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_control_slave_write),      //                          .write
		.ctrl_writedata       (mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_control_slave_writedata),  //                          .writedata
		.ctrl_readdata        (mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_control_slave_readdata),   //                          .readdata
		.buf_byteenable       (mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_buffer_slave_byteenable),  //  avalon_char_buffer_slave.byteenable
		.buf_chipselect       (mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_buffer_slave_chipselect),  //                          .chipselect
		.buf_read             (mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_buffer_slave_read),        //                          .read
		.buf_write            (mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_buffer_slave_write),       //                          .write
		.buf_writedata        (mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_buffer_slave_writedata),   //                          .writedata
		.buf_readdata         (mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_buffer_slave_readdata),    //                          .readdata
		.buf_waitrequest      (mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_buffer_slave_waitrequest), //                          .waitrequest
		.buf_address          (mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_buffer_slave_address),     //                          .address
		.stream_ready         (video_character_buffer_with_dma_0_avalon_char_source_ready),                               //        avalon_char_source.ready
		.stream_startofpacket (video_character_buffer_with_dma_0_avalon_char_source_startofpacket),                       //                          .startofpacket
		.stream_endofpacket   (video_character_buffer_with_dma_0_avalon_char_source_endofpacket),                         //                          .endofpacket
		.stream_valid         (video_character_buffer_with_dma_0_avalon_char_source_valid),                               //                          .valid
		.stream_data          (video_character_buffer_with_dma_0_avalon_char_source_data)                                 //                          .data
	);

	MMIX_system_video_dual_clock_buffer_0 video_dual_clock_buffer_0 (
		.clk_stream_in            (clocks_sys_clk_clk),                                                 //         clock_stream_in.clk
		.reset_stream_in          (rst_controller_reset_out_reset),                                     //   clock_stream_in_reset.reset
		.clk_stream_out           (video_pll_0_vga_clk_clk),                                            //        clock_stream_out.clk
		.reset_stream_out         (rst_controller_002_reset_out_reset),                                 //  clock_stream_out_reset.reset
		.stream_in_ready          (video_character_buffer_with_dma_0_avalon_char_source_ready),         //   avalon_dc_buffer_sink.ready
		.stream_in_startofpacket  (video_character_buffer_with_dma_0_avalon_char_source_startofpacket), //                        .startofpacket
		.stream_in_endofpacket    (video_character_buffer_with_dma_0_avalon_char_source_endofpacket),   //                        .endofpacket
		.stream_in_valid          (video_character_buffer_with_dma_0_avalon_char_source_valid),         //                        .valid
		.stream_in_data           (video_character_buffer_with_dma_0_avalon_char_source_data),          //                        .data
		.stream_out_ready         (video_dual_clock_buffer_0_avalon_dc_buffer_source_ready),            // avalon_dc_buffer_source.ready
		.stream_out_startofpacket (video_dual_clock_buffer_0_avalon_dc_buffer_source_startofpacket),    //                        .startofpacket
		.stream_out_endofpacket   (video_dual_clock_buffer_0_avalon_dc_buffer_source_endofpacket),      //                        .endofpacket
		.stream_out_valid         (video_dual_clock_buffer_0_avalon_dc_buffer_source_valid),            //                        .valid
		.stream_out_data          (video_dual_clock_buffer_0_avalon_dc_buffer_source_data)              //                        .data
	);

	MMIX_system_video_vga_controller_0 video_vga_controller_0 (
		.clk           (video_pll_0_vga_clk_clk),                                         //        clock_reset.clk
		.reset         (rst_controller_002_reset_out_reset),                              //  clock_reset_reset.reset
		.data          (video_dual_clock_buffer_0_avalon_dc_buffer_source_data),          //    avalon_vga_sink.data
		.startofpacket (video_dual_clock_buffer_0_avalon_dc_buffer_source_startofpacket), //                   .startofpacket
		.endofpacket   (video_dual_clock_buffer_0_avalon_dc_buffer_source_endofpacket),   //                   .endofpacket
		.valid         (video_dual_clock_buffer_0_avalon_dc_buffer_source_valid),         //                   .valid
		.ready         (video_dual_clock_buffer_0_avalon_dc_buffer_source_ready),         //                   .ready
		.VGA_CLK       (vga_wire_CLK),                                                    // external_interface.export
		.VGA_HS        (vga_wire_HS),                                                     //                   .export
		.VGA_VS        (vga_wire_VS),                                                     //                   .export
		.VGA_R         (vga_wire_R),                                                      //                   .export
		.VGA_G         (vga_wire_G),                                                      //                   .export
		.VGA_B         (vga_wire_B)                                                       //                   .export
	);

	MMIX_system_video_pll_0 video_pll_0 (
		.ref_clk_clk        (clocks_sys_clk_clk),             //      ref_clk.clk
		.ref_reset_reset    (rst_controller_reset_out_reset), //    ref_reset.reset
		.vga_clk_clk        (video_pll_0_vga_clk_clk),        //      vga_clk.clk
		.reset_source_reset (video_pll_0_reset_source_reset)  // reset_source.reset
	);

	MMIX_system_mm_interconnect_0 mm_interconnect_0 (
		.clocks_sys_clk_clk                                                                (clocks_sys_clk_clk),                                                                                  //                                                        clocks_sys_clk.clk
		.mmix_qsys_0_reset_n_reset_bridge_in_reset_reset                                   (rst_controller_reset_out_reset),                                                                      //                             mmix_qsys_0_reset_n_reset_bridge_in_reset.reset
		.sdram_reset_reset_bridge_in_reset_reset                                           (rst_controller_reset_out_reset),                                                                      //                                     sdram_reset_reset_bridge_in_reset.reset
		.mmix_qsys_0_master_address                                                        (mmix_qsys_0_master_address),                                                                          //                                                    mmix_qsys_0_master.address
		.mmix_qsys_0_master_waitrequest                                                    (mmix_qsys_0_master_waitrequest),                                                                      //                                                                      .waitrequest
		.mmix_qsys_0_master_byteenable                                                     (mmix_qsys_0_master_byteenable),                                                                       //                                                                      .byteenable
		.mmix_qsys_0_master_read                                                           (mmix_qsys_0_master_read),                                                                             //                                                                      .read
		.mmix_qsys_0_master_readdata                                                       (mmix_qsys_0_master_readdata),                                                                         //                                                                      .readdata
		.mmix_qsys_0_master_readdatavalid                                                  (mmix_qsys_0_master_readdatavalid),                                                                    //                                                                      .readdatavalid
		.mmix_qsys_0_master_write                                                          (mmix_qsys_0_master_write),                                                                            //                                                                      .write
		.mmix_qsys_0_master_writedata                                                      (mmix_qsys_0_master_writedata),                                                                        //                                                                      .writedata
		.Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_data_address              (mm_interconnect_0_altera_up_flash_memory_ip_core_avalon_interface_0_flash_data_address),              //          Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_data.address
		.Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_data_write                (mm_interconnect_0_altera_up_flash_memory_ip_core_avalon_interface_0_flash_data_write),                //                                                                      .write
		.Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_data_read                 (mm_interconnect_0_altera_up_flash_memory_ip_core_avalon_interface_0_flash_data_read),                 //                                                                      .read
		.Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_data_readdata             (mm_interconnect_0_altera_up_flash_memory_ip_core_avalon_interface_0_flash_data_readdata),             //                                                                      .readdata
		.Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_data_writedata            (mm_interconnect_0_altera_up_flash_memory_ip_core_avalon_interface_0_flash_data_writedata),            //                                                                      .writedata
		.Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_data_byteenable           (mm_interconnect_0_altera_up_flash_memory_ip_core_avalon_interface_0_flash_data_byteenable),           //                                                                      .byteenable
		.Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_data_waitrequest          (mm_interconnect_0_altera_up_flash_memory_ip_core_avalon_interface_0_flash_data_waitrequest),          //                                                                      .waitrequest
		.Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_data_chipselect           (mm_interconnect_0_altera_up_flash_memory_ip_core_avalon_interface_0_flash_data_chipselect),           //                                                                      .chipselect
		.Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_erase_control_write       (mm_interconnect_0_altera_up_flash_memory_ip_core_avalon_interface_0_flash_erase_control_write),       // Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_erase_control.write
		.Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_erase_control_read        (mm_interconnect_0_altera_up_flash_memory_ip_core_avalon_interface_0_flash_erase_control_read),        //                                                                      .read
		.Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_erase_control_readdata    (mm_interconnect_0_altera_up_flash_memory_ip_core_avalon_interface_0_flash_erase_control_readdata),    //                                                                      .readdata
		.Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_erase_control_writedata   (mm_interconnect_0_altera_up_flash_memory_ip_core_avalon_interface_0_flash_erase_control_writedata),   //                                                                      .writedata
		.Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_erase_control_byteenable  (mm_interconnect_0_altera_up_flash_memory_ip_core_avalon_interface_0_flash_erase_control_byteenable),  //                                                                      .byteenable
		.Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_erase_control_waitrequest (mm_interconnect_0_altera_up_flash_memory_ip_core_avalon_interface_0_flash_erase_control_waitrequest), //                                                                      .waitrequest
		.Altera_UP_Flash_Memory_IP_Core_Avalon_Interface_0_flash_erase_control_chipselect  (mm_interconnect_0_altera_up_flash_memory_ip_core_avalon_interface_0_flash_erase_control_chipselect),  //                                                                      .chipselect
		.sdram_s1_address                                                                  (mm_interconnect_0_sdram_s1_address),                                                                  //                                                              sdram_s1.address
		.sdram_s1_write                                                                    (mm_interconnect_0_sdram_s1_write),                                                                    //                                                                      .write
		.sdram_s1_read                                                                     (mm_interconnect_0_sdram_s1_read),                                                                     //                                                                      .read
		.sdram_s1_readdata                                                                 (mm_interconnect_0_sdram_s1_readdata),                                                                 //                                                                      .readdata
		.sdram_s1_writedata                                                                (mm_interconnect_0_sdram_s1_writedata),                                                                //                                                                      .writedata
		.sdram_s1_byteenable                                                               (mm_interconnect_0_sdram_s1_byteenable),                                                               //                                                                      .byteenable
		.sdram_s1_readdatavalid                                                            (mm_interconnect_0_sdram_s1_readdatavalid),                                                            //                                                                      .readdatavalid
		.sdram_s1_waitrequest                                                              (mm_interconnect_0_sdram_s1_waitrequest),                                                              //                                                                      .waitrequest
		.sdram_s1_chipselect                                                               (mm_interconnect_0_sdram_s1_chipselect),                                                               //                                                                      .chipselect
		.video_character_buffer_with_dma_0_avalon_char_buffer_slave_address                (mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_buffer_slave_address),                //            video_character_buffer_with_dma_0_avalon_char_buffer_slave.address
		.video_character_buffer_with_dma_0_avalon_char_buffer_slave_write                  (mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_buffer_slave_write),                  //                                                                      .write
		.video_character_buffer_with_dma_0_avalon_char_buffer_slave_read                   (mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_buffer_slave_read),                   //                                                                      .read
		.video_character_buffer_with_dma_0_avalon_char_buffer_slave_readdata               (mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_buffer_slave_readdata),               //                                                                      .readdata
		.video_character_buffer_with_dma_0_avalon_char_buffer_slave_writedata              (mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_buffer_slave_writedata),              //                                                                      .writedata
		.video_character_buffer_with_dma_0_avalon_char_buffer_slave_byteenable             (mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_buffer_slave_byteenable),             //                                                                      .byteenable
		.video_character_buffer_with_dma_0_avalon_char_buffer_slave_waitrequest            (mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_buffer_slave_waitrequest),            //                                                                      .waitrequest
		.video_character_buffer_with_dma_0_avalon_char_buffer_slave_chipselect             (mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_buffer_slave_chipselect),             //                                                                      .chipselect
		.video_character_buffer_with_dma_0_avalon_char_control_slave_address               (mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_control_slave_address),               //           video_character_buffer_with_dma_0_avalon_char_control_slave.address
		.video_character_buffer_with_dma_0_avalon_char_control_slave_write                 (mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_control_slave_write),                 //                                                                      .write
		.video_character_buffer_with_dma_0_avalon_char_control_slave_read                  (mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_control_slave_read),                  //                                                                      .read
		.video_character_buffer_with_dma_0_avalon_char_control_slave_readdata              (mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_control_slave_readdata),              //                                                                      .readdata
		.video_character_buffer_with_dma_0_avalon_char_control_slave_writedata             (mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_control_slave_writedata),             //                                                                      .writedata
		.video_character_buffer_with_dma_0_avalon_char_control_slave_byteenable            (mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_control_slave_byteenable),            //                                                                      .byteenable
		.video_character_buffer_with_dma_0_avalon_char_control_slave_chipselect            (mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_control_slave_chipselect)             //                                                                      .chipselect
	);

	MMIX_system_irq_mapper irq_mapper (
		.clk        (),                      //       clk.clk
		.reset      (),                      // clk_reset.reset
		.sender_irq (mmix_qsys_0_d_irq_irq)  //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                 // reset_in0.reset
		.clk            (clocks_sys_clk_clk),             //       clk.clk
		.reset_out      (rst_controller_reset_out_reset), // reset_out.reset
		.reset_req      (),                               // (terminated)
		.reset_req_in0  (1'b0),                           // (terminated)
		.reset_in1      (1'b0),                           // (terminated)
		.reset_req_in1  (1'b0),                           // (terminated)
		.reset_in2      (1'b0),                           // (terminated)
		.reset_req_in2  (1'b0),                           // (terminated)
		.reset_in3      (1'b0),                           // (terminated)
		.reset_req_in3  (1'b0),                           // (terminated)
		.reset_in4      (1'b0),                           // (terminated)
		.reset_req_in4  (1'b0),                           // (terminated)
		.reset_in5      (1'b0),                           // (terminated)
		.reset_req_in5  (1'b0),                           // (terminated)
		.reset_in6      (1'b0),                           // (terminated)
		.reset_req_in6  (1'b0),                           // (terminated)
		.reset_in7      (1'b0),                           // (terminated)
		.reset_req_in7  (1'b0),                           // (terminated)
		.reset_in8      (1'b0),                           // (terminated)
		.reset_req_in8  (1'b0),                           // (terminated)
		.reset_in9      (1'b0),                           // (terminated)
		.reset_req_in9  (1'b0),                           // (terminated)
		.reset_in10     (1'b0),                           // (terminated)
		.reset_req_in10 (1'b0),                           // (terminated)
		.reset_in11     (1'b0),                           // (terminated)
		.reset_req_in11 (1'b0),                           // (terminated)
		.reset_in12     (1'b0),                           // (terminated)
		.reset_req_in12 (1'b0),                           // (terminated)
		.reset_in13     (1'b0),                           // (terminated)
		.reset_req_in13 (1'b0),                           // (terminated)
		.reset_in14     (1'b0),                           // (terminated)
		.reset_req_in14 (1'b0),                           // (terminated)
		.reset_in15     (1'b0),                           // (terminated)
		.reset_req_in15 (1'b0)                            // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.clk            (clk_clk),                            //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_002 (
		.reset_in0      (video_pll_0_reset_source_reset),     // reset_in0.reset
		.clk            (video_pll_0_vga_clk_clk),            //       clk.clk
		.reset_out      (rst_controller_002_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
